module vsync()
//1920x1080 lab monitors


endmodule